module univeral(
  
